/*
 --------------------------------------------------------------------------
   Pegasus - Copyright (C) 2012 Gregory Matthew James.

   This file is part of Pegasus.

   Pegasus is free; you can redistribute it and/or modify
   it under the terms of the GNU General Public License as published by
   the Free Software Foundation; either version 3 of the License, or
   (at your option) any later version.

   Pegasus is distributed in the hope that it will be useful,
   but WITHOUT ANY WARRANTY; without even the implied warranty of
   MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE. See the
   GNU General Public License for more details.

   You should have received a copy of the GNU General Public License
   along with this program. If not, see <http://www.gnu.org/licenses/>.
 --------------------------------------------------------------------------
*/

/*
 --------------------------------------------------------------------------
 -- Project Code      : pegasus
 -- Interface Name    : clk_rst_sync_intf
 -- Author            : mammenx
 -- Function          : This interface encapsulates a typical clock & its
                        associated synchronous reset signal.
 --------------------------------------------------------------------------
*/

interface clk_rst_sync_intf  (input logic clk_ir,  rst_sync_l);

  //Modport
  modport sync  (
                  input clk_ir, rst_sync_l
                );

endinterface  //  clk_rst_sync_intf

/*
 --------------------------------------------------------------------------

 -- <Header>
 

 -- <Log>

[08-06-2014  02:25:23 PM][mammenx] Moved under intf directory

[08-06-2014  02:20:11 PM][mammenx] Initial Commit

[28-05-14 20:18:21] [mammenx] Moved log section to bottom of file

 --------------------------------------------------------------------------
*/
